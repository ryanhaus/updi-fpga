// testbench 
