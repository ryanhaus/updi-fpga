module top (
	input clk,
	input rst,
	input start,
	output updi
);

	// 

endmodule
