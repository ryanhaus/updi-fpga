enum {
	UPDI_LDS,
	UPDI_LD,
	UPDI_STS,
	UPDI_ST,
	UPDI_LDCS,
	UPDI_REPEAT,
	UPDI_STCS,
	UPDI_KEY
} updi_instruction;

module updi_interface (

);

endmodule
