// Module for handling UART TX traffic
/* verilator lint_off WIDTHEXPAND */
module uart_tx #(
	parameter DATA_BITS = 8, // 5 - 9
	parameter PARITY_BIT = "none", // "none", "even", or "odd"
	parameter STOP_BITS = 1 // 1 - 2
) (
	input clk, // baud rate for UART
	input rst,

	input [DATA_BITS-1 : 0] tx_data,
	input start,
	output logic ready,
	output logic tx
);

	uart_state state;
	logic [DATA_BITS-1 : 0] data;
	logic [$clog2(DATA_BITS)-1 : 0] counter; // used for data & stop bits

	// parity module
	logic parity_result;
	parity #(.BITS(DATA_BITS)) parity_inst (data, parity_result);

	// UART state machine
	always_ff @(posedge clk) begin
		if (rst) begin
			state = UART_IDLE;
			ready = 'b0;
			tx = 'b1;
		end
		else begin
			case (state)
				UART_IDLE: begin
					// idle is 1
					ready = 'b1;
					tx = 'b1;

					// handle going to start bit
					if (start) begin
						state = UART_START;
						ready = 'b0;
						data = tx_data;
						counter = 'b0;
					end
				end

				UART_START: begin
					// always one 0 bit
					tx = 'b0;
					state = UART_DATA;
				end

				UART_DATA: begin
					// handle transmission
					tx = data[counter]; // LSB

					// handle going to next state if applicable
					if (counter == DATA_BITS-1) begin
						counter = 'b0;

						if (PARITY_BIT == "none") begin
							state = UART_STOP;
						end
						else begin
							state = UART_PARITY;
						end
					end
					else begin
						// otherwise just keep going through data bits
						counter = counter + 'b1;
						state = UART_DATA;
					end
				end

				UART_PARITY: begin
					// handle parity, parity_result is always odd parity
					case (PARITY_BIT)
						"even": tx = ~parity_result;
						"odd": tx = parity_result;
					endcase

					state = UART_STOP;
				end

				UART_STOP: begin
					// handle stop bit(s)
					tx = 'b1;

					counter = counter + 'b1;
					if (counter < STOP_BITS) begin
						// have to repeat for multiple stop bits
						state = UART_STOP;
					end
					else begin
						// handle next state
						// TODO: for speed, skip going back to IDLE if start is 1
						state = UART_IDLE;
						ready = 'b1;
					end
				end
			endcase
		end
	end

endmodule
/* lint_on */
